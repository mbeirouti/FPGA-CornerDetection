library IEEE;

use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use std.textio.all;

entity squares is
	

	port(
		clk : in std_logic;
		xGrad : in std_logic_vector(7 downto 0);
		yGrad : in std_logic_vector(7 downto 0);
		xGradSq : out std_logic_vector(15 downto 0);
		yGradSq: out std_logic_vector(15 downto 0);
		xyGrad : out std_logic_vector(15 downto 0));

end squares;


architecture implementation of squares is
	
	
	
	begin


	
	
	
	


end implementation;