library IEEE;

use ieee.std_logic_1164.all;

entity PixelManagementUnit_tb is
end entity;

architecture PixelManagementUnit_tst of PixelManagementUnit_tb is

begin

end architecture;