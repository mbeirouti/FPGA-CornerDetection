library IEEE;

entity TriIntMemory is

	port (
		yIn, xIn, xyIn: in integer;
		yOut,xOut,xyOut: out integer
	);
	
end entity;

architecture TriIntMemory_Impl of TriIntMemory is

begin

end architecture;